module BigAlu(ai,bi,Aluop2,Aluop,ri);
input Aluop2;
wire MSB_wire,lessi;
wire [31:0] cci;
wire V;
input [2:0] Aluop;
input [31:0] ai;
input [31:0] bi;
output Z;
wire Z1,elde;
output [31:0] ri;
Alu1 th1(ai[0],bi[0],Aluop2,Aluop2,MSB_wire,Aluop[0],Aluop[1],cci[1],ri[0]);
Alu1 th2(ai[1],bi[1],cci[1],Aluop[2],1'b0,Aluop[0],Aluop[1],cci[2],ri[1]);
Alu1 th3(ai[2],bi[2],cci[2],Aluop[2],1'b0,Aluop[0],Aluop[1],cci[3],ri[2]);
Alu1 th4(ai[3],bi[3],cci[3],Aluop[2],1'b0,Aluop[0],Aluop[1],cci[4],ri[3]);
Alu1 th5(ai[4],bi[4],cci[4],Aluop[2],1'b0,Aluop[0],Aluop[1],cci[5],ri[4]);
Alu1 th6(ai[5],bi[5],cci[5],Aluop[2],1'b0,Aluop[0],Aluop[1],cci[6],ri[5]);
Alu1 th7(ai[6],bi[6],cci[6],Aluop[2],1'b0,Aluop[0],Aluop[1],cci[7],ri[6]);
Alu1 th8(ai[7],bi[7],cci[7],Aluop[2],1'b0,Aluop[0],Aluop[1],cci[8],ri[7]);
Alu1 th9(ai[8],bi[8],cci[8],Aluop[2],1'b0,Aluop[0],Aluop[1],cci[9],ri[8]);
Alu1 th10(ai[9],bi[9],cci[9],Aluop[2],1'b0,Aluop[0],Aluop[1],cci[10],ri[9]);
Alu1 th11(ai[10],bi[10],cci[10],Aluop[2],1'b0,Aluop[0],Aluop[1],cci[11],ri[10]);
Alu1 th12(ai[11],bi[11],cci[11],Aluop[2],1'b0,Aluop[0],Aluop[1],cci[12],ri[11]);
Alu1 th13(ai[12],bi[12],cci[12],Aluop[2],1'b0,Aluop[0],Aluop[1],cci[13],ri[12]);
Alu1 th14(ai[13],bi[13],cci[13],Aluop[2],1'b0,Aluop[0],Aluop[1],cci[14],ri[13]);
Alu1 th15(ai[14],bi[14],cci[14],Aluop[2],1'b0,Aluop[0],Aluop[1],cci[15],ri[14]);
Alu1 th16(ai[15],bi[15],cci[15],Aluop[2],1'b0,Aluop[0],Aluop[1],cci[16],ri[15]);
Alu1 th17(ai[16],bi[16],cci[16],Aluop[2],1'b0,Aluop[0],Aluop[1],cci[17],ri[16]);
Alu1 th18(ai[17],bi[17],cci[17],Aluop[2],1'b0,Aluop[0],Aluop[1],cci[18],ri[17]);
Alu1 th119(ai[18],bi[18],cci[18],Aluop[2],1'b0,Aluop[0],Aluop[1],cci[19],ri[18]);
Alu1 th20(ai[19],bi[19],cci[19],Aluop[2],1'b0,Aluop[0],Aluop[1],cci[20],ri[19]);
Alu1 th21(ai[20],bi[20],cci[20],Aluop[2],1'b0,Aluop[0],Aluop[1],cci[21],ri[20]);
Alu1 th22(ai[21],bi[21],cci[21],Aluop[2],1'b0,Aluop[0],Aluop[1],cci[22],ri[21]);
Alu1 th23(ai[22],bi[22],cci[22],Aluop[2],1'b0,Aluop[0],Aluop[1],cci[23],ri[22]);
Alu1 th24(ai[23],bi[23],cci[23],Aluop[2],1'b0,Aluop[0],Aluop[1],cci[24],ri[23]);
Alu1 th25(ai[24],bi[24],cci[24],Aluop[2],1'b0,Aluop[0],Aluop[1],cci[25],ri[24]);
Alu1 th26(ai[25],bi[25],cci[25],Aluop[2],1'b0,Aluop[0],Aluop[1],cci[26],ri[25]);
Alu1 th27(ai[26],bi[26],cci[26],Aluop[2],1'b0,Aluop[0],Aluop[1],cci[27],ri[26]);
Alu1 th28(ai[27],bi[27],cci[27],Aluop[2],1'b0,Aluop[0],Aluop[1],cci[28],ri[27]);
Alu1 th29(ai[28],bi[28],cci[28],Aluop[2],1'b0,Aluop[0],Aluop[1],cci[29],ri[28]);
Alu1 th30(ai[29],bi[29],cci[29],Aluop[2],1'b0,Aluop[0],Aluop[1],cci[30],ri[29]);
Alu1 th31(ai[30],bi[30],cci[30],Aluop[2],1'b0,Aluop[0],Aluop[1],cci[31],ri[30]);
MSBALU alu(ai[31],bi[31],cci[31],Aluop[0],Aluop[1],Aluop[2],1'b0,ri[31],MSB_wire,elde,V);
or orsonuc(Z1,ri[0],ri[1],ri[2],ri[3],ri[4],ri[5],ri[6],ri[7],ri[8],ri[9],ri[10],ri[11],ri[12],ri[13],ri[14],ri[15],ri[16],ri[17],ri[18],ri[19],ri[20],ri[21],ri[22],ri[23],ri[24],ri[25],ri[26],ri[27],ri[28],ri[29],ri[30],ri[31]);
not notsonuc(Z,Z1);
endmodule